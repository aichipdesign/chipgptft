4. Executing CHECK pass (checking for obvious problems).
Checking module Decoder...
Found and reported 0 problems.

End of script. Logfile hash: 9504430b16, CPU: user 0.01s system 0.00s, MEM: 11.37 MB peak
